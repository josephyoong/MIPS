// sign_extend
// Sign Extend

module sign_extend #(
) (
    input [15:0] I;
    output [31:0] O;
);

endmodule
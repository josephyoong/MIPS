// PC_plus4
// PC Plus 4

module PC_plus4 #(
) (
    input [31:0] I;
    output [31:0] O;
);

assign O = I + 4;

endmodule
// PC
// Program Counter (PC)

module PC #(
) (
    input clk,
    input [31:0] PC_next,
    output [31:0] PC
);

endmodule
// data_memory
// Data Memory

module data_memory #(
) (
    input clk,
    input WE; // write enable
    input [31:0] WD, // write data
    input [31:0] A,
    output [31:0] RD,
);

endmodule
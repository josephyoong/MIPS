// PC_branch
// Program Counter (PC) Branch 

module PC_branch (
) (
    input [31:0] I;
    
);

endmodule
// instruction_memory
// Instruction Memory

module instruction_memory #(
) (
    input clk,
    input [31:0] A,
    output [31:0] RD,
);

endmodule